interface Mem;
endinterface

(* synthesize *)
module mkMem(Mem);
endmodule: mkMem
