import Mem::*;

(* synthesize *)
module mkTop(Empty);
    Mem mem <- mkMem;
endmodule: mkTop